`ifndef HLX_INTFC_SVH
`define HLX_INTFC_SVH

`define AXI_MM_AW 64
`define AXI_MM_DW 512
`define AXI_LITE_AW 32
`define AXI_LITE_DW 32


`endif /* HLX_INTFC_SVH */
