// Sanjay Rai (sanjay.d.rai@gmail.com)
//
`timescale 1 ps / 1 ps

module shell_top (
  inout [3:0]BMC_GPIO_tri_io,
  input BMC_UART_rxd,
  output BMC_UART_txd,
  input C1_SYS_CLK_clk_n,
  input C1_SYS_CLK_clk_p,
  input [7:0]C0_DDR_SREF_CTRL_IN,
  output [7:0]C0_DDR_SREF_CTRL_OUT,
  input [7:0]C2_DDR_SREF_CTRL_IN,
  output [7:0]C2_DDR_SREF_CTRL_OUT,
  input [7:0]C3_DDR_SREF_CTRL_IN,
  output [7:0]C3_DDR_SREF_CTRL_OUT,
  hlx_AXI_LITE_intfc.master M_AXI_LITE_TO_HLS_PR_NORTH, 
  hlx_AXI_MM_intfc.slave S_AXI_MM_MIG, 
  hlx_AXI_MM_intfc.slave S_AXI_MM_PCIM, 
  output axi_reset_n_out,
  output c1_ddr4_act_n,
  output [16:0]c1_ddr4_adr,
  output [1:0]c1_ddr4_ba,
  output [1:0]c1_ddr4_bg,
  output [0:0]c1_ddr4_ck_c,
  output [0:0]c1_ddr4_ck_t,
  output [0:0]c1_ddr4_cke,
  output [0:0]c1_ddr4_cs_n,
  inout [71:0]c1_ddr4_dq,
  inout [17:0]c1_ddr4_dqs_c,
  inout [17:0]c1_ddr4_dqs_t,
  output [0:0]c1_ddr4_odt,
  output c1_ddr4_par,
  output c1_ddr4_reset_n,
  output c1_init_calib_complete,
  output clk_out_125M,
  output clk_out_300M,
  output clk_out_400M,
  output clk_out_250M,
  output clk_out_PROG,
  inout iic_scl_io,
  inout iic_sda_io,
  input [15:0]pcie_mgt_rxn,
  input [15:0]pcie_mgt_rxp,
  output [15:0]pcie_mgt_txn,
  output [15:0]pcie_mgt_txp,
  output rst_main_n,
  output MIG_0_RST_N,
  output MIG_2_RST_N,
  output MIG_3_RST_N,
  output RESET_GATE,
  input sys_clk,
  input sys_clk_gt,
  input sys_rst_n);

  wire [3:0]BMC_GPIO_tri_i;
  wire [3:0]BMC_GPIO_tri_io;
  wire [3:0]BMC_GPIO_tri_o;
  wire [3:0]BMC_GPIO_tri_t;

  wire iic_scl_i;
  wire iic_scl_o;
  wire iic_scl_t;
  wire iic_sda_i;
  wire iic_sda_o;
  wire iic_sda_t;



  PCIe_Bridge_ICAP_complex PCIe_Bridge_ICAP_complex_i (
        .BMC_GPIO_tri_i(BMC_GPIO_tri_i),
        .BMC_GPIO_tri_o(BMC_GPIO_tri_o),
        .BMC_GPIO_tri_t(BMC_GPIO_tri_t),
        .BMC_UART_rxd(BMC_UART_rxd),
        .BMC_UART_txd(BMC_UART_txd),
        .C1_SYS_CLK_clk_n(C1_SYS_CLK_clk_n),
        .C1_SYS_CLK_clk_p(C1_SYS_CLK_clk_p),
        .C0_DDR_SREF_CTRL_IN(C0_DDR_SREF_CTRL_IN),
        .C0_DDR_SREF_CTRL_OUT(C0_DDR_SREF_CTRL_OUT),
        .C2_DDR_SREF_CTRL_IN(C2_DDR_SREF_CTRL_IN),
        .C2_DDR_SREF_CTRL_OUT(C2_DDR_SREF_CTRL_OUT),
        .C3_DDR_SREF_CTRL_IN(C3_DDR_SREF_CTRL_IN),
        .C3_DDR_SREF_CTRL_OUT(C3_DDR_SREF_CTRL_OUT),
        .MIG_0_RST_N(MIG_0_RST_N),
        .MIG_2_RST_N(MIG_2_RST_N),
        .MIG_3_RST_N(MIG_3_RST_N),
        .M_AXI_LITE_TO_HLS_PR_NORTH_araddr(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_araddr),
        .M_AXI_LITE_TO_HLS_PR_NORTH_arprot(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_arprot),
        .M_AXI_LITE_TO_HLS_PR_NORTH_arready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_arready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_arvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_arvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awaddr(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awaddr),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awprot(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awprot),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_awvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_awvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_bready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_bready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_bresp(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_bresp),
        .M_AXI_LITE_TO_HLS_PR_NORTH_bvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_bvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rdata(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rdata),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rresp(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rresp),
        .M_AXI_LITE_TO_HLS_PR_NORTH_rvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_rvalid),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wdata(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wdata),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wready(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wready),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wstrb(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wstrb),
        .M_AXI_LITE_TO_HLS_PR_NORTH_wvalid(M_AXI_LITE_TO_HLS_PR_NORTH.AXI_LITE_wvalid),
        .RESET_GATE(RESET_GATE),
        .S_AXI_MM_0_araddr(S_AXI_MM_MIG.AXI_araddr),
        .S_AXI_MM_0_arburst(S_AXI_MM_MIG.AXI_arburst),
        .S_AXI_MM_0_arcache(S_AXI_MM_MIG.AXI_arcache),
        .S_AXI_MM_0_arid(S_AXI_MM_MIG.AXI_arid),
        .S_AXI_MM_0_arlen(S_AXI_MM_MIG.AXI_arlen),
        .S_AXI_MM_0_arlock(S_AXI_MM_MIG.AXI_arlock),
        .S_AXI_MM_0_arprot(S_AXI_MM_MIG.AXI_arprot),
        .S_AXI_MM_0_arqos(S_AXI_MM_MIG.AXI_arqos),
        .S_AXI_MM_0_arready(S_AXI_MM_MIG.AXI_arready),
        .S_AXI_MM_0_arregion(S_AXI_MM_MIG.AXI_arregion),
        .S_AXI_MM_0_arsize(S_AXI_MM_MIG.AXI_arsize),
        .S_AXI_MM_0_arvalid(S_AXI_MM_MIG.AXI_arvalid),
        .S_AXI_MM_0_awaddr(S_AXI_MM_MIG.AXI_awaddr),
        .S_AXI_MM_0_awburst(S_AXI_MM_MIG.AXI_awburst),
        .S_AXI_MM_0_awcache(S_AXI_MM_MIG.AXI_awcache),
        .S_AXI_MM_0_awid(S_AXI_MM_MIG.AXI_awid),
        .S_AXI_MM_0_awlen(S_AXI_MM_MIG.AXI_awlen),
        .S_AXI_MM_0_awlock(S_AXI_MM_MIG.AXI_awlock),
        .S_AXI_MM_0_awprot(S_AXI_MM_MIG.AXI_awprot),
        .S_AXI_MM_0_awqos(S_AXI_MM_MIG.AXI_awqos),
        .S_AXI_MM_0_awready(S_AXI_MM_MIG.AXI_awready),
        .S_AXI_MM_0_awregion(S_AXI_MM_MIG.AXI_awregion),
        .S_AXI_MM_0_awsize(S_AXI_MM_MIG.AXI_awsize),
        .S_AXI_MM_0_awvalid(S_AXI_MM_MIG.AXI_awvalid),
        .S_AXI_MM_0_bid(S_AXI_MM_MIG.AXI_bid),
        .S_AXI_MM_0_bready(S_AXI_MM_MIG.AXI_bready),
        .S_AXI_MM_0_bresp(S_AXI_MM_MIG.AXI_bresp),
        .S_AXI_MM_0_bvalid(S_AXI_MM_MIG.AXI_bvalid),
        .S_AXI_MM_0_rdata(S_AXI_MM_MIG.AXI_rdata),
        .S_AXI_MM_0_rid(S_AXI_MM_MIG.AXI_rid),
        .S_AXI_MM_0_rlast(S_AXI_MM_MIG.AXI_rlast),
        .S_AXI_MM_0_rready(S_AXI_MM_MIG.AXI_rready),
        .S_AXI_MM_0_rresp(S_AXI_MM_MIG.AXI_rresp),
        .S_AXI_MM_0_rvalid(S_AXI_MM_MIG.AXI_rvalid),
        .S_AXI_MM_0_wdata(S_AXI_MM_MIG.AXI_wdata),
        .S_AXI_MM_0_wlast(S_AXI_MM_MIG.AXI_wlast),
        .S_AXI_MM_0_wready(S_AXI_MM_MIG.AXI_wready),
        .S_AXI_MM_0_wstrb(S_AXI_MM_MIG.AXI_wstrb),
        .S_AXI_MM_0_wvalid(S_AXI_MM_MIG.AXI_wvalid),
        .S_AXI_MM_PCIM_araddr(S_AXI_MM_PCIM.AXI_araddr),
        .S_AXI_MM_PCIM_arburst(S_AXI_MM_PCIM.AXI_arburst),
        .S_AXI_MM_PCIM_arcache(S_AXI_MM_PCIM.AXI_arcache),
        .S_AXI_MM_PCIM_arid(S_AXI_MM_PCIM.AXI_arid),
        .S_AXI_MM_PCIM_arlen(S_AXI_MM_PCIM.AXI_arlen),
        .S_AXI_MM_PCIM_arlock(S_AXI_MM_PCIM.AXI_arlock),
        .S_AXI_MM_PCIM_arprot(S_AXI_MM_PCIM.AXI_arprot),
        .S_AXI_MM_PCIM_arqos(S_AXI_MM_PCIM.AXI_arqos),
        .S_AXI_MM_PCIM_arready(S_AXI_MM_PCIM.AXI_arready),
        .S_AXI_MM_PCIM_arregion(S_AXI_MM_PCIM.AXI_arregion),
        .S_AXI_MM_PCIM_arsize(S_AXI_MM_PCIM.AXI_arsize),
        .S_AXI_MM_PCIM_arvalid(S_AXI_MM_PCIM.AXI_arvalid),
        .S_AXI_MM_PCIM_awaddr(S_AXI_MM_PCIM.AXI_awaddr),
        .S_AXI_MM_PCIM_awburst(S_AXI_MM_PCIM.AXI_awburst),
        .S_AXI_MM_PCIM_awcache(S_AXI_MM_PCIM.AXI_awcache),
        .S_AXI_MM_PCIM_awid(S_AXI_MM_PCIM.AXI_awid),
        .S_AXI_MM_PCIM_awlen(S_AXI_MM_PCIM.AXI_awlen),
        .S_AXI_MM_PCIM_awlock(S_AXI_MM_PCIM.AXI_awlock),
        .S_AXI_MM_PCIM_awprot(S_AXI_MM_PCIM.AXI_awprot),
        .S_AXI_MM_PCIM_awqos(S_AXI_MM_PCIM.AXI_awqos),
        .S_AXI_MM_PCIM_awready(S_AXI_MM_PCIM.AXI_awready),
        .S_AXI_MM_PCIM_awregion(S_AXI_MM_PCIM.AXI_awregion),
        .S_AXI_MM_PCIM_awsize(S_AXI_MM_PCIM.AXI_awsize),
        .S_AXI_MM_PCIM_awvalid(S_AXI_MM_PCIM.AXI_awvalid),
        .S_AXI_MM_PCIM_bid(S_AXI_MM_PCIM.AXI_bid),
        .S_AXI_MM_PCIM_bready(S_AXI_MM_PCIM.AXI_bready),
        .S_AXI_MM_PCIM_bresp(S_AXI_MM_PCIM.AXI_bresp),
        .S_AXI_MM_PCIM_bvalid(S_AXI_MM_PCIM.AXI_bvalid),
        .S_AXI_MM_PCIM_rdata(S_AXI_MM_PCIM.AXI_rdata),
        .S_AXI_MM_PCIM_rid(S_AXI_MM_PCIM.AXI_rid),
        .S_AXI_MM_PCIM_rlast(S_AXI_MM_PCIM.AXI_rlast),
        .S_AXI_MM_PCIM_rready(S_AXI_MM_PCIM.AXI_rready),
        .S_AXI_MM_PCIM_rresp(S_AXI_MM_PCIM.AXI_rresp),
        .S_AXI_MM_PCIM_rvalid(S_AXI_MM_PCIM.AXI_rvalid),
        .S_AXI_MM_PCIM_wdata(S_AXI_MM_PCIM.AXI_wdata),
        .S_AXI_MM_PCIM_wlast(S_AXI_MM_PCIM.AXI_wlast),
        .S_AXI_MM_PCIM_wready(S_AXI_MM_PCIM.AXI_wready),
        .S_AXI_MM_PCIM_wstrb(S_AXI_MM_PCIM.AXI_wstrb),
        .S_AXI_MM_PCIM_wvalid(S_AXI_MM_PCIM.AXI_wvalid),
        .axi_reset_n_250M_out(axi_reset_n_out),
        .c1_ddr4_act_n(c1_ddr4_act_n),
        .c1_ddr4_adr(c1_ddr4_adr),
        .c1_ddr4_ba(c1_ddr4_ba),
        .c1_ddr4_bg(c1_ddr4_bg),
        .c1_ddr4_ck_c(c1_ddr4_ck_c),
        .c1_ddr4_ck_t(c1_ddr4_ck_t),
        .c1_ddr4_cke(c1_ddr4_cke),
        .c1_ddr4_cs_n(c1_ddr4_cs_n),
        .c1_ddr4_par(c1_ddr4_par),
        .c1_ddr4_dq(c1_ddr4_dq),
        .c1_ddr4_dqs_c(c1_ddr4_dqs_c),
        .c1_ddr4_dqs_t(c1_ddr4_dqs_t),
        .c1_ddr4_odt(c1_ddr4_odt),
        .c1_ddr4_reset_n(c1_ddr4_reset_n),
        .c1_init_calib_complete(c1_init_calib_complete),
        .clk_out_125M(clk_out_125M),
        .clk_out_250M(clk_out_250M),
        .clk_out_300M(clk_out_300M),
        .clk_out_400M(clk_out_400M),
        .clk_out_PROG(clk_out_PROG),
        .iic_scl_i(iic_scl_i),
        .iic_scl_o(iic_scl_o),
        .iic_scl_t(iic_scl_t),
        .iic_sda_i(iic_sda_i),
        .iic_sda_o(iic_sda_o),
        .iic_sda_t(iic_sda_t),
        .pcie_mgt_rxn(pcie_mgt_rxn),
        .pcie_mgt_rxp(pcie_mgt_rxp),
        .pcie_mgt_txn(pcie_mgt_txn),
        .pcie_mgt_txp(pcie_mgt_txp),
        .rst_main_n(rst_main_n),
        .sys_clk(sys_clk),
        .sys_clk_gt(sys_clk_gt),
        .sys_rst_n(sys_rst_n));

  IOBUF iic_scl_iobuf
       (.I(iic_scl_o),
        .IO(iic_scl_io),
        .O(iic_scl_i),
        .T(iic_scl_t));
  IOBUF iic_sda_iobuf
       (.I(iic_sda_o),
        .IO(iic_sda_io),
        .O(iic_sda_i),
        .T(iic_sda_t));

  genvar i;
  generate
    for (i=0; i < 4; i++) begin
      IOBUF BMC_GPIO_tri_iobuf
           (.I(BMC_GPIO_tri_o[i]),
            .IO(BMC_GPIO_tri_io[i]),
            .O(BMC_GPIO_tri_i[i]),
            .T(BMC_GPIO_tri_t[i]));
    end
  endgenerate

endmodule
